`define IMPORT_HOSTIF 
`define XILINX_SYS_CLK 
`define DataBusWidth 256
`define USE_WIDE_WIDTH 
`define ConnectalVersion 18.08.1
`define NumberOfMasters 1
`define PinType Top_Pins
`define PinTypeInclude FlashTop
`define NumberOfUserTiles 1
`define SlaveDataBusWidth 32
`define SlaveControlAddrWidth 5
`define BurstLenSize 10
`define project_dir $(DTOP)
`define MainClockPeriod 8
`define DerivedClockPeriod 9.091000
`define PcieClockPeriod 4
`define XILINX 1
`define VirtexUltrascale 
`define XilinxUltrascale 
`define PCIE 
`define PCIE3 
`define PcieHostInterface 
`define PhysAddrWidth 40
`define NUMBER_OF_LEDS 2
`define PcieLanes 8
`define CONNECTAL_BITS_DEPENDENCES hw/mkTop.bit
`define CONNECTAL_RUN_SCRIPT $(CONNECTALDIR)/scripts/run.pcietest
`define BOARD_vcu108 
