
#include "GeneratedTypes.h"


