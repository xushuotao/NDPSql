typedef enum{Byte, Short, Int, Long, BigInt} SimdMode deriving (Bits, Eq, FShow); //3-bit
